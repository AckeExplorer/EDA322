use library